library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

use work.Types.all;

entity tb is 
end entity;

architecture beh of tb is
begin
end architecture beh;
